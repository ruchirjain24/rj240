//https://drive.google.com/file/d/1axWmpz-saQrbXKGRZL8bU9B34uWZ7vvR/view
module hello;
 initial
 begin
 $display("Hello World");
 $finish ;
 end
endmodule